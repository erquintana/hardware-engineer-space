module tb
    always @() // always_comb, always_ff, always_latch
endmodule