class driver();
    
endclass