//------------------------------------------------------------------------------
// Project: Verifying the VeriRISC CPU
// File:    veriRISC_CPU.sv
// Author:  Esteban Rodríguez Quintana
// Date:    <>
//
// Description: <>
//
// Revision History:
// - <Date>: <Version / Modification Description>
//
//------------------------------------------------------------------------------

