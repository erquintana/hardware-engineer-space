`include "universal_reg.sv"

module tb;

    
endmodule