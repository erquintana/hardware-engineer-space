module fifo(
    input clock, rd_en, wr_en, rst_n, 
    input [7:0] data_in;
    output full, empty,
    output reg [7:0] data_out
);


endmodule